module controls(
  output reg [7:0] vol1, //Information about relative volume
  output reg [7:0] vol2,
  output reg [7:0] vol3,
  output reg [7:0] vol4,
  output reg [7:0] freq1, //Information about frequency, may not literally be frequency
  output reg [7:0] freq2,
  output reg [7:0] freq3,
  output reg [7:0] freq4
);
  //And then actually make the module
endmodule
