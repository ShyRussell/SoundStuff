// Sabrina Pereira, Shy Russell, Jonah Spicher
/*-----------------------------------------------------------------------------
Square Wave Generator
-----------------------------------------------------------------------------*/
`include "register.v"
`include "counter.v"

module square_wave
#(parameter resolution_bits = 8, parameter counter_width = 8)
(
    output [resolution_bits-1:0] square_out,
    input  clk,   // System clock
    input  [counter_width-1:0] frequency_control  // Control for the output frequency

);

// Wires for D-flip-flop that generates square wave
wire  [resolution_bits-1:0]  d_to_q_inv; // Wire ~q to d
reg  inv_trigger; //Tell when to invert signal

// Wires for counter MAY NEED TO BE LARGER
wire  [counter_width-1:0]  count;


d_flip_flop sqwave_generator(.q(square_out),.q_inv(d_to_q_inv),.d(d_to_q_inv),.clk(inv_trigger));

counter counter(.count(count),.clk(clk),.reset(inv_trigger));


// Controls for reset and waves
always @* begin
if (count == frequency_control)
  inv_trigger=1;
else
  inv_trigger=0;
end

always @(frequency_control) begin
  inv_trigger=1;
end

endmodule

module sound_square_wave
#(parameter resolution_bits = 8, parameter counter_width = 8)
(
    output reg [resolution_bits-1:0] square_out,
    input  clk,   // System clock
    input  [counter_width-1:0] frequency_control  // Control for the output frequency

);

// Wires for D-flip-flop that generates square wave
wire  [resolution_bits-2:0]  d_to_q_inv, sq_wave; // Wire ~q to d
reg  inv_trigger; //Tell when to invert signal

// Wires for counter MAY NEED TO BE LARGER
wire  [counter_width-1:0]  count;

d_flip_flop #(7) sqwave_generator(.q(sq_wave),.q_inv(d_to_q_inv),.d(d_to_q_inv),.clk(inv_trigger));

counter counter(.count(count),.clk(clk),.reset(inv_trigger));



// Controls for reset and waves
always @* begin
square_out = {!sq_wave[0], sq_wave};
if (count == frequency_control)
  inv_trigger=1;
else
  inv_trigger=0;
end

always @(frequency_control) begin
  inv_trigger=1;
end

endmodule
